// 512-point Real-valued FFT Engine (via 256-point complex FFT)
// Exploits conjugate symmetry of real inputs: packs 512 real samples into 256
// complex values, runs a standard radix-2 DIT FFT, then unscrambles the result
// to recover 256 unique frequency bins.
//
// Data flow: COLLECT 512 real samples (packed pairwise into 256 complex)
//          → COMPUTE 8 butterfly stages (standard 256-point complex FFT)
//          → UNSCRAMBLE + magnitude output (256 bins)
//
// Uses Q1.14 fixed-point twiddle factors loaded from twiddle.hex.
// The twiddle ROM stores W_512^k for k=0..255 (256 entries).
// Butterfly stages access at even addresses: W_256^k = W_512^(2k).
//
// Memory: same 2× DP16KD as a 256-point complex FFT (no increase).
// Requires twiddle.hex with 256 entries (generated by gen_twiddle.py).

module fft_real512 (
    input  wire        clk,
    input  wire        rst_n,

    // Input sample stream (real-valued, 16-bit signed)
    input  wire signed [15:0] sample_in,
    input  wire               sample_valid,

    // Output magnitude (sequential during output phase)
    output reg  [7:0]  mag_addr,
    output reg  [8:0]  mag_data,
    output reg         mag_valid,

    // Status
    output wire        busy
);

    // ======================================================================
    // Constants
    // ======================================================================
    localparam N = 256;  // Complex FFT size (processes 2*N real samples)

    // FSM states
    localparam [1:0] S_COLLECT    = 2'd0,
                     S_COMPUTE    = 2'd1,
                     S_UNSCRAMBLE = 2'd2;

    reg [1:0] state;
    assign busy = (state != S_COLLECT);

    // ======================================================================
    // Dual-port RAM for real and imaginary parts
    // Two always blocks per array = true dual-port → ECP5 DP16KD inference
    // ======================================================================
    (* no_rw_check *) reg [15:0] re_mem [0:N-1];
    (* no_rw_check *) reg [15:0] im_mem [0:N-1];

    // Port A and B control signals (directly driven by combinational mux)
    reg [7:0]  re_addr_a, re_addr_b;
    reg [15:0] re_wdata_a, re_wdata_b;
    reg        re_we_a, re_we_b;
    reg [7:0]  im_addr_a, im_addr_b;
    reg [15:0] im_wdata_a, im_wdata_b;
    reg        im_we_a, im_we_b;

    // Registered read outputs (1-cycle latency)
    reg [15:0] re_rdata_a, re_rdata_b;
    reg [15:0] im_rdata_a, im_rdata_b;

    // Real part: port A
    always @(posedge clk) begin
        if (re_we_a) re_mem[re_addr_a] <= re_wdata_a;
        re_rdata_a <= re_mem[re_addr_a];
    end
    // Real part: port B
    always @(posedge clk) begin
        if (re_we_b) re_mem[re_addr_b] <= re_wdata_b;
        re_rdata_b <= re_mem[re_addr_b];
    end
    // Imaginary part: port A
    always @(posedge clk) begin
        if (im_we_a) im_mem[im_addr_a] <= im_wdata_a;
        im_rdata_a <= im_mem[im_addr_a];
    end
    // Imaginary part: port B
    always @(posedge clk) begin
        if (im_we_b) im_mem[im_addr_b] <= im_wdata_b;
        im_rdata_b <= im_mem[im_addr_b];
    end

    // ======================================================================
    // Twiddle factor ROM: 256 entries x 32 bits {cos[15:0], sin[15:0]}
    // Q1.14 format (scale = 16384), registered read for block ROM inference
    // Stores W_512^k for k=0..255.
    // Butterfly uses W_256^j = W_512^(2j) → address = 2*j.
    // Unscramble uses W_512^k directly → address = k.
    // ======================================================================
    reg [31:0] twiddle [0:N-1];
    initial $readmemh("twiddle.hex", twiddle);

    reg [7:0]  tw_addr;
    reg [31:0] tw_rdata;
    always @(posedge clk) tw_rdata <= twiddle[tw_addr];

    // ======================================================================
    // Bit-reverse function for DIT input reordering (8-bit for N=256)
    // ======================================================================
    function [7:0] bit_reverse;
        input [7:0] idx;
        bit_reverse = {idx[0], idx[1], idx[2], idx[3],
                       idx[4], idx[5], idx[6], idx[7]};
    endfunction

    // ======================================================================
    // Collection counter and sample pairing register
    // ======================================================================
    reg [8:0] sample_count;           // 0..511 (9-bit)
    reg signed [15:0] even_sample;    // Holds x[2n] while waiting for x[2n+1]

    // ======================================================================
    // Butterfly state
    // ======================================================================
    reg [2:0] bfly_stage;    // FFT stage (0..7)
    reg [6:0] bfly_idx;      // Butterfly index within stage (0..127)
    reg [1:0] bfly_step;     // Sub-step within butterfly (0..2)

    // ======================================================================
    // Butterfly address computation
    // Insert a 0/1 at bit position 'bfly_stage' to get addresses p and q
    // ======================================================================
    reg [7:0] addr_p_calc, addr_q_calc;
    reg [6:0] tw_addr_calc;

    always @(*) begin
        case (bfly_stage)
            3'd0: begin
                addr_p_calc  = {bfly_idx, 1'b0};
                addr_q_calc  = {bfly_idx, 1'b1};
                tw_addr_calc = 7'd0;
            end
            3'd1: begin
                addr_p_calc  = {bfly_idx[6:1], 1'b0, bfly_idx[0]};
                addr_q_calc  = {bfly_idx[6:1], 1'b1, bfly_idx[0]};
                tw_addr_calc = {bfly_idx[0], 6'd0};
            end
            3'd2: begin
                addr_p_calc  = {bfly_idx[6:2], 1'b0, bfly_idx[1:0]};
                addr_q_calc  = {bfly_idx[6:2], 1'b1, bfly_idx[1:0]};
                tw_addr_calc = {bfly_idx[1:0], 5'd0};
            end
            3'd3: begin
                addr_p_calc  = {bfly_idx[6:3], 1'b0, bfly_idx[2:0]};
                addr_q_calc  = {bfly_idx[6:3], 1'b1, bfly_idx[2:0]};
                tw_addr_calc = {bfly_idx[2:0], 4'd0};
            end
            3'd4: begin
                addr_p_calc  = {bfly_idx[6:4], 1'b0, bfly_idx[3:0]};
                addr_q_calc  = {bfly_idx[6:4], 1'b1, bfly_idx[3:0]};
                tw_addr_calc = {bfly_idx[3:0], 3'd0};
            end
            3'd5: begin
                addr_p_calc  = {bfly_idx[6:5], 1'b0, bfly_idx[4:0]};
                addr_q_calc  = {bfly_idx[6:5], 1'b1, bfly_idx[4:0]};
                tw_addr_calc = {bfly_idx[4:0], 2'd0};
            end
            3'd6: begin
                addr_p_calc  = {bfly_idx[6], 1'b0, bfly_idx[5:0]};
                addr_q_calc  = {bfly_idx[6], 1'b1, bfly_idx[5:0]};
                tw_addr_calc = {bfly_idx[5:0], 1'd0};
            end
            3'd7: begin
                addr_p_calc  = {1'b0, bfly_idx[6:0]};
                addr_q_calc  = {1'b1, bfly_idx[6:0]};
                tw_addr_calc = bfly_idx[6:0];
            end
        endcase
    end

    // ======================================================================
    // Butterfly computation pipeline
    // ======================================================================

    // Latched values from registered RAM reads
    reg signed [15:0] a_re, a_im;
    reg signed [15:0] b_re, b_im;
    reg signed [15:0] tw_cos_r, tw_sin_r;
    reg [7:0] addr_p_r, addr_q_r;

    // Complex twiddle multiply: W * B
    // W = cos - j*sin, so W*B = (cos*Bre + sin*Bim) + j(cos*Bim - sin*Bre)
    /* verilator lint_off UNUSEDSIGNAL */
    wire signed [31:0] tw_x_re = tw_cos_r * b_re + tw_sin_r * b_im;
    wire signed [31:0] tw_x_im = tw_cos_r * b_im - tw_sin_r * b_re;
    /* verilator lint_on UNUSEDSIGNAL */

    // Scale twiddle product back from Q1.14 (arithmetic right shift by 14)
    wire signed [17:0] t_re = tw_x_re[31:14];
    wire signed [17:0] t_im = tw_x_im[31:14];

    // Butterfly results with 1/2 scaling per stage
    wire signed [17:0] a_re_ext = {{2{a_re[15]}}, a_re};
    wire signed [17:0] a_im_ext = {{2{a_im[15]}}, a_im};

    /* verilator lint_off UNUSEDSIGNAL */
    wire signed [17:0] sum_re = a_re_ext + t_re;
    wire signed [17:0] sum_im = a_im_ext + t_im;
    wire signed [17:0] dif_re = a_re_ext - t_re;
    wire signed [17:0] dif_im = a_im_ext - t_im;
    /* verilator lint_on UNUSEDSIGNAL */

    // Arithmetic right shift by 1, truncate to 16 bits
    wire [15:0] p_re_new = sum_re[16:1];
    wire [15:0] p_im_new = sum_im[16:1];
    wire [15:0] q_re_new = dif_re[16:1];
    wire [15:0] q_im_new = dif_im[16:1];

    // ======================================================================
    // Unscramble state
    // ======================================================================
    reg [7:0] unscr_k;       // Current output bin index (0..255)
    reg [1:0] unscr_step;    // Pipeline sub-step (0..2)
    reg [7:0] unscr_k_d;     // Delayed k for output alignment

    // Unscramble registered intermediate values
    // Ze[k] = (Z[k] + Z*[(N-k)%N]) / 2
    // Zo[k] = (Z[k] - Z*[(N-k)%N]) / (2j)
    //
    // In component form (Zm = Z[(N-k)%N]):
    //   Ze_re = (Zk_re + Zm_re) / 2     Ze_im = (Zk_im - Zm_im) / 2
    //   Zo_re = (Zk_im + Zm_im) / 2     Zo_im = (Zm_re - Zk_re) / 2
    //
    // We register the half-scaled values to keep 16-bit width for the
    // twiddle multiply (matching the butterfly's 16x16 multiplier structure).
    reg signed [15:0] ze_re_r, ze_im_r;
    reg signed [15:0] zo_re_r, zo_im_r;

    // Unscramble twiddle multiply: W_512^k * Zo[k]
    // Reuses the same structure as the butterfly: cos*re + sin*im, cos*im - sin*re
    // tw_cos_r and tw_sin_r are loaded in unscr_step 1.
    // zo_re_r and zo_im_r are loaded in unscr_step 1.
    /* verilator lint_off UNUSEDSIGNAL */
    wire signed [31:0] wzo_re = tw_cos_r * zo_re_r + tw_sin_r * zo_im_r;
    wire signed [31:0] wzo_im = tw_cos_r * zo_im_r - tw_sin_r * zo_re_r;
    /* verilator lint_on UNUSEDSIGNAL */

    // X[k] = Ze[k] + W_512^k * Zo[k]
    // Ze values are already /2 scaled (16-bit).
    // W*Zo product needs >>14 for Q1.14 de-scaling.
    wire signed [17:0] ze_re_ext = {{2{ze_re_r[15]}}, ze_re_r};
    wire signed [17:0] ze_im_ext = {{2{ze_im_r[15]}}, ze_im_r};
    wire signed [17:0] wzo_re_s  = wzo_re[31:14];
    wire signed [17:0] wzo_im_s  = wzo_im[31:14];

    /* verilator lint_off UNUSEDSIGNAL */
    wire signed [17:0] x_re_full = ze_re_ext + wzo_re_s;
    wire signed [17:0] x_im_full = ze_im_ext + wzo_im_s;
    /* verilator lint_on UNUSEDSIGNAL */

    // ======================================================================
    // Magnitude computation (used during UNSCRAMBLE phase)
    // ======================================================================
    // Take upper 16 bits of the 18-bit X values (discard 2 LSBs for magnitude)
    wire signed [15:0] x_re_mag = x_re_full[17:2];
    wire signed [15:0] x_im_mag = x_im_full[17:2];

    wire [15:0] abs_re = x_re_mag[15] ? (~x_re_mag + 16'd1) : x_re_mag;
    wire [15:0] abs_im = x_im_mag[15] ? (~x_im_mag + 16'd1) : x_im_mag;
    wire [15:0] mag_max = (abs_re > abs_im) ? abs_re : abs_im;
    /* verilator lint_off UNUSEDSIGNAL */
    wire [15:0] mag_min = (abs_re > abs_im) ? abs_im : abs_re;
    /* verilator lint_on UNUSEDSIGNAL */
    // Approximate magnitude: max + min/4 (within ~5% of true magnitude)
    wire [15:0] magnitude = mag_max + {2'b00, mag_min[15:2]};

    // Log2 magnitude via priority encoder (4.4 fixed-point)
    // Gives ~96 dB dynamic range mapped to 0-440 pixel range
    reg [3:0] log2_int;
    /* verilator lint_off UNUSEDSIGNAL */
    reg [15:0] mag_norm;
    /* verilator lint_on UNUSEDSIGNAL */
    always @(*) begin
        log2_int = 4'd0;
        mag_norm = 16'd0;
        if      (magnitude[15]) begin log2_int = 4'd15; mag_norm = magnitude;        end
        else if (magnitude[14]) begin log2_int = 4'd14; mag_norm = magnitude << 1;   end
        else if (magnitude[13]) begin log2_int = 4'd13; mag_norm = magnitude << 2;   end
        else if (magnitude[12]) begin log2_int = 4'd12; mag_norm = magnitude << 3;   end
        else if (magnitude[11]) begin log2_int = 4'd11; mag_norm = magnitude << 4;   end
        else if (magnitude[10]) begin log2_int = 4'd10; mag_norm = magnitude << 5;   end
        else if (magnitude[9])  begin log2_int = 4'd9;  mag_norm = magnitude << 6;   end
        else if (magnitude[8])  begin log2_int = 4'd8;  mag_norm = magnitude << 7;   end
        else if (magnitude[7])  begin log2_int = 4'd7;  mag_norm = magnitude << 8;   end
        else if (magnitude[6])  begin log2_int = 4'd6;  mag_norm = magnitude << 9;   end
        else if (magnitude[5])  begin log2_int = 4'd5;  mag_norm = magnitude << 10;  end
        else if (magnitude[4])  begin log2_int = 4'd4;  mag_norm = magnitude << 11;  end
        else if (magnitude[3])  begin log2_int = 4'd3;  mag_norm = magnitude << 12;  end
        else if (magnitude[2])  begin log2_int = 4'd2;  mag_norm = magnitude << 13;  end
        else if (magnitude[1])  begin log2_int = 4'd1;  mag_norm = magnitude << 14;  end
        else if (magnitude[0])  begin log2_int = 4'd0;  mag_norm = 16'h8000;         end
    end
    wire [3:0] log2_frac = mag_norm[14:11];
    wire [7:0] log2_val  = {log2_int, log2_frac};
    // Scale 4.4 fixed-point log2 (0-255) to 0-438 pixel range: (val * 440) >> 8
    /* verilator lint_off UNUSEDSIGNAL */
    wire [16:0] log2_scaled = log2_val * 9'd440;
    /* verilator lint_on UNUSEDSIGNAL */
    wire [8:0]  capped_mag = (magnitude == 16'd0) ? 9'd0 : log2_scaled[16:8];

    // ======================================================================
    // RAM port address/control mux (directly drives dual-port RAM signals)
    // ======================================================================
    always @(*) begin
        // Defaults: no writes, address 0
        re_addr_a  = 8'd0;  re_addr_b  = 8'd0;
        re_wdata_a = 16'd0; re_wdata_b = 16'd0;
        re_we_a    = 1'b0;  re_we_b    = 1'b0;
        im_addr_a  = 8'd0;  im_addr_b  = 8'd0;
        im_wdata_a = 16'd0; im_wdata_b = 16'd0;
        im_we_a    = 1'b0;  im_we_b    = 1'b0;
        tw_addr    = 8'd0;

        case (state)
            S_COLLECT: begin
                // Write paired samples on odd counts:
                // re_mem[bit_rev(n)] = even_sample, im_mem[bit_rev(n)] = sample_in
                re_addr_a  = bit_reverse(sample_count[8:1]);
                re_wdata_a = even_sample;
                re_we_a    = sample_valid & sample_count[0];
                im_addr_a  = bit_reverse(sample_count[8:1]);
                im_wdata_a = sample_in;
                im_we_a    = sample_valid & sample_count[0];
            end

            S_COMPUTE: begin
                // Butterfly twiddle: W_256^j = W_512^(2j)
                tw_addr = {tw_addr_calc, 1'b0};
                case (bfly_step)
                    2'd0: begin
                        // Read setup: present addresses for registered read
                        re_addr_a = addr_p_calc;
                        re_addr_b = addr_q_calc;
                        im_addr_a = addr_p_calc;
                        im_addr_b = addr_q_calc;
                    end
                    2'd1: begin
                        // Read data is now available in rdata registers
                        // (latching into a_re/b_re happens in state machine)
                    end
                    2'd2: begin
                        // Write butterfly results via both ports
                        re_addr_a  = addr_p_r;
                        re_addr_b  = addr_q_r;
                        re_wdata_a = p_re_new;
                        re_wdata_b = q_re_new;
                        re_we_a    = 1'b1;
                        re_we_b    = 1'b1;
                        im_addr_a  = addr_p_r;
                        im_addr_b  = addr_q_r;
                        im_wdata_a = p_im_new;
                        im_wdata_b = q_im_new;
                        im_we_a    = 1'b1;
                        im_we_b    = 1'b1;
                    end
                    default: ;
                endcase
            end

            S_UNSCRAMBLE: begin
                // Read Z[k] from port A, Z[(N-k)%N] from port B
                re_addr_a = unscr_k;
                im_addr_a = unscr_k;
                re_addr_b = (unscr_k == 8'd0) ? 8'd0 : (8'd0 - unscr_k);
                im_addr_b = (unscr_k == 8'd0) ? 8'd0 : (8'd0 - unscr_k);
                // Twiddle for unscramble: W_512^k, addressed directly
                tw_addr   = unscr_k;
            end

            default: ;
        endcase
    end

    // ======================================================================
    // Main state machine
    // ======================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state        <= S_COLLECT;
            sample_count <= 9'd0;
            even_sample  <= 16'd0;
            bfly_stage   <= 3'd0;
            bfly_idx     <= 7'd0;
            bfly_step    <= 2'd0;
            unscr_k      <= 8'd0;
            unscr_step   <= 2'd0;
            unscr_k_d    <= 8'd0;
            mag_valid    <= 1'b0;
            mag_addr     <= 8'd0;
            mag_data     <= 9'd0;
            ze_re_r      <= 16'd0;
            ze_im_r      <= 16'd0;
            zo_re_r      <= 16'd0;
            zo_im_r      <= 16'd0;
            a_re         <= 16'd0;
            a_im         <= 16'd0;
            b_re         <= 16'd0;
            b_im         <= 16'd0;
            tw_cos_r     <= 16'd0;
            tw_sin_r     <= 16'd0;
            addr_p_r     <= 8'd0;
            addr_q_r     <= 8'd0;
        end else begin
            mag_valid <= 1'b0;  // Default: no output

            case (state)
                // ----------------------------------------------------------
                // COLLECT: Store 512 real samples, packed pairwise as complex.
                // Even samples (count[0]==0) are latched in even_sample.
                // Odd samples (count[0]==1) trigger a write:
                //   re_mem[bit_rev(n)] = even_sample (x[2n])
                //   im_mem[bit_rev(n)] = sample_in   (x[2n+1])
                // Writes are driven by the combinational mux above.
                // ----------------------------------------------------------
                S_COLLECT: begin
                    if (sample_valid) begin
                        if (!sample_count[0]) begin
                            // Even sample: latch and wait for odd partner
                            even_sample <= sample_in;
                        end
                        // Odd sample: write is handled by combinational mux

                        if (sample_count == 9'd511) begin
                            sample_count <= 9'd0;
                            bfly_stage   <= 3'd0;
                            bfly_idx     <= 7'd0;
                            bfly_step    <= 2'd0;
                            state        <= S_COMPUTE;
                        end else begin
                            sample_count <= sample_count + 9'd1;
                        end
                    end
                end

                // ----------------------------------------------------------
                // COMPUTE: 8 stages x 128 butterflies x 3 cycles each
                // (Identical to fft256 except twiddle address doubled in mux)
                // Step 0: present addresses (RAM reads on next posedge)
                // Step 1: latch registered read data + twiddle
                // Step 2: write butterfly results (via mux), advance
                // ----------------------------------------------------------
                S_COMPUTE: begin
                    case (bfly_step)
                        2'd0: begin
                            // Addresses driven by mux; latch for write-back
                            addr_p_r  <= addr_p_calc;
                            addr_q_r  <= addr_q_calc;
                            bfly_step <= 2'd1;
                        end
                        2'd1: begin
                            // Registered reads are now valid; latch into butterfly regs
                            a_re     <= $signed(re_rdata_a);
                            a_im     <= $signed(im_rdata_a);
                            b_re     <= $signed(re_rdata_b);
                            b_im     <= $signed(im_rdata_b);
                            tw_cos_r <= $signed(tw_rdata[31:16]);
                            tw_sin_r <= $signed(tw_rdata[15:0]);
                            bfly_step <= 2'd2;
                        end
                        2'd2: begin
                            // Writes driven by mux; advance to next butterfly
                            bfly_step <= 2'd0;
                            if (bfly_idx == 7'd127) begin
                                bfly_idx <= 7'd0;
                                if (bfly_stage == 3'd7) begin
                                    unscr_k    <= 8'd0;
                                    unscr_step <= 2'd0;
                                    state      <= S_UNSCRAMBLE;
                                end else begin
                                    bfly_stage <= bfly_stage + 3'd1;
                                end
                            end else begin
                                bfly_idx <= bfly_idx + 7'd1;
                            end
                        end
                        default: bfly_step <= 2'd0;
                    endcase
                end

                // ----------------------------------------------------------
                // UNSCRAMBLE: Recover 512-point real FFT bins from 256-point
                // complex FFT results, then compute log2 magnitude.
                //
                // For bin k (0..255):
                //   Z[k]  from port A,  Z[(N-k)%N] from port B
                //   Ze[k] = (Z[k] + Z*[(N-k)%N]) / 2
                //   Zo[k] = (Z[k] - Z*[(N-k)%N]) / (2j)
                //   X[k]  = Ze[k] + W_512^k * Zo[k]
                //
                // Step 0: present addresses (RAM/ROM reads on next posedge)
                // Step 1: latch data, compute Ze and Zo
                // Step 2: magnitude of X[k] → output
                // ----------------------------------------------------------
                S_UNSCRAMBLE: begin
                    case (unscr_step)
                        2'd0: begin
                            // Addresses driven by mux; save k for output
                            unscr_k_d  <= unscr_k;
                            unscr_step <= 2'd1;
                        end
                        2'd1: begin
                            // RAM/ROM data valid. Compute Ze and Zo components.
                            // Zk = (re_rdata_a, im_rdata_a)
                            // Zm = (re_rdata_b, im_rdata_b) = Z[(N-k)%N]
                            // Z*m = (Zm_re, -Zm_im)
                            //
                            // Ze = (Zk + Z*m) / 2:
                            //   Ze_re = (Zk_re + Zm_re) >>> 1
                            //   Ze_im = (Zk_im - Zm_im) >>> 1
                            //
                            // Zo = (Zk - Z*m) / (2j) = -j*(Zk - Z*m) / 2:
                            //   Zo_re = (Zk_im + Zm_im) >>> 1
                            //   Zo_im = (Zm_re - Zk_re) >>> 1
                            ze_re_r <= ($signed(re_rdata_a) + $signed(re_rdata_b)) >>> 1;
                            ze_im_r <= ($signed(im_rdata_a) - $signed(im_rdata_b)) >>> 1;
                            zo_re_r <= ($signed(im_rdata_a) + $signed(im_rdata_b)) >>> 1;
                            zo_im_r <= ($signed(re_rdata_b) - $signed(re_rdata_a)) >>> 1;

                            // Latch twiddle W_512^k
                            tw_cos_r <= $signed(tw_rdata[31:16]);
                            tw_sin_r <= $signed(tw_rdata[15:0]);

                            unscr_step <= 2'd2;
                        end
                        2'd2: begin
                            // Multiply + magnitude computed combinationally above.
                            // Output the result.
                            mag_addr  <= unscr_k_d;
                            mag_data  <= capped_mag;
                            mag_valid <= 1'b1;
                            unscr_step <= 2'd0;
                            if (unscr_k == 8'd255) begin
                                unscr_k <= 8'd0;
                                state   <= S_COLLECT;
                            end else begin
                                unscr_k <= unscr_k + 8'd1;
                            end
                        end
                        default: unscr_step <= 2'd0;
                    endcase
                end

                default: state <= S_COLLECT;
            endcase
        end
    end

endmodule
