// 256-point Radix-2 DIT FFT Engine
// Accepts 16-bit signed samples one at a time, computes in-place FFT,
// and outputs magnitude values suitable for spectrum display.
//
// Data flow: COLLECT 256 samples → COMPUTE 8 butterfly stages → MAGNITUDE → output
// Uses Q1.14 fixed-point twiddle factors loaded from twiddle.hex.
// Each butterfly stage scales by 1/2 to prevent overflow (total 1/N normalization).
//
// Memory is structured as dual-port RAM for ECP5 block RAM (EBR) inference.
// Requires twiddle.hex in the working directory (generated by gen_twiddle.py).

module fft256 #(
    parameter MAG_SHIFT = 3   // Right-shift magnitude before capping at display range
) (
    input  wire        clk,
    input  wire        rst_n,

    // Input sample stream
    input  wire signed [15:0] sample_in,
    input  wire               sample_valid,

    // Output magnitude (sequential during output phase)
    output reg  [7:0]  mag_addr,
    output reg  [8:0]  mag_data,
    output reg         mag_valid,

    // Status
    output wire        busy
);

    // ======================================================================
    // Constants
    // ======================================================================
    localparam N      = 256;
    localparam LOG2_N = 8;
    localparam [8:0] MAX_MAG = 9'd440;

    // FSM states
    localparam [1:0] S_COLLECT   = 2'd0,
                     S_COMPUTE   = 2'd1,
                     S_MAGNITUDE = 2'd2;

    reg [1:0] state;
    assign busy = (state != S_COLLECT);

    // ======================================================================
    // Dual-port RAM for real and imaginary parts
    // Two always blocks per array = true dual-port → ECP5 DP16KD inference
    // ======================================================================
    (* no_rw_check *) reg [15:0] re_mem [0:N-1];
    (* no_rw_check *) reg [15:0] im_mem [0:N-1];

    // Port A and B control signals (directly driven by combinational mux)
    reg [7:0]  re_addr_a, re_addr_b;
    reg [15:0] re_wdata_a, re_wdata_b;
    reg        re_we_a, re_we_b;
    reg [7:0]  im_addr_a, im_addr_b;
    reg [15:0] im_wdata_a, im_wdata_b;
    reg        im_we_a, im_we_b;

    // Registered read outputs (1-cycle latency)
    reg [15:0] re_rdata_a, re_rdata_b;
    reg [15:0] im_rdata_a, im_rdata_b;

    // Real part: port A
    always @(posedge clk) begin
        if (re_we_a) re_mem[re_addr_a] <= re_wdata_a;
        re_rdata_a <= re_mem[re_addr_a];
    end
    // Real part: port B
    always @(posedge clk) begin
        if (re_we_b) re_mem[re_addr_b] <= re_wdata_b;
        re_rdata_b <= re_mem[re_addr_b];
    end
    // Imaginary part: port A
    always @(posedge clk) begin
        if (im_we_a) im_mem[im_addr_a] <= im_wdata_a;
        im_rdata_a <= im_mem[im_addr_a];
    end
    // Imaginary part: port B
    always @(posedge clk) begin
        if (im_we_b) im_mem[im_addr_b] <= im_wdata_b;
        im_rdata_b <= im_mem[im_addr_b];
    end

    // ======================================================================
    // Twiddle factor ROM: 128 entries x 32 bits {cos[15:0], sin[15:0]}
    // Q1.14 format (scale = 16384), registered read for block ROM inference
    // ======================================================================
    reg [31:0] twiddle [0:127];
    initial $readmemh("twiddle.hex", twiddle);

    reg [6:0]  tw_addr;
    reg [31:0] tw_rdata;
    always @(posedge clk) tw_rdata <= twiddle[tw_addr];

    // ======================================================================
    // Bit-reverse function for DIT input reordering
    // ======================================================================
    function [7:0] bit_reverse;
        input [7:0] idx;
        bit_reverse = {idx[0], idx[1], idx[2], idx[3],
                       idx[4], idx[5], idx[6], idx[7]};
    endfunction

    // ======================================================================
    // Collection counter
    // ======================================================================
    reg [7:0] sample_count;

    // ======================================================================
    // Butterfly state
    // ======================================================================
    reg [2:0] bfly_stage;    // FFT stage (0..7)
    reg [6:0] bfly_idx;      // Butterfly index within stage (0..127)
    reg [1:0] bfly_step;     // Sub-step within butterfly (0..2)

    // ======================================================================
    // Butterfly address computation
    // Insert a 0/1 at bit position 'bfly_stage' to get addresses p and q
    // ======================================================================
    reg [7:0] addr_p_calc, addr_q_calc;
    reg [6:0] tw_addr_calc;

    always @(*) begin
        case (bfly_stage)
            3'd0: begin
                addr_p_calc  = {bfly_idx, 1'b0};
                addr_q_calc  = {bfly_idx, 1'b1};
                tw_addr_calc = 7'd0;
            end
            3'd1: begin
                addr_p_calc  = {bfly_idx[6:1], 1'b0, bfly_idx[0]};
                addr_q_calc  = {bfly_idx[6:1], 1'b1, bfly_idx[0]};
                tw_addr_calc = {bfly_idx[0], 6'd0};
            end
            3'd2: begin
                addr_p_calc  = {bfly_idx[6:2], 1'b0, bfly_idx[1:0]};
                addr_q_calc  = {bfly_idx[6:2], 1'b1, bfly_idx[1:0]};
                tw_addr_calc = {bfly_idx[1:0], 5'd0};
            end
            3'd3: begin
                addr_p_calc  = {bfly_idx[6:3], 1'b0, bfly_idx[2:0]};
                addr_q_calc  = {bfly_idx[6:3], 1'b1, bfly_idx[2:0]};
                tw_addr_calc = {bfly_idx[2:0], 4'd0};
            end
            3'd4: begin
                addr_p_calc  = {bfly_idx[6:4], 1'b0, bfly_idx[3:0]};
                addr_q_calc  = {bfly_idx[6:4], 1'b1, bfly_idx[3:0]};
                tw_addr_calc = {bfly_idx[3:0], 3'd0};
            end
            3'd5: begin
                addr_p_calc  = {bfly_idx[6:5], 1'b0, bfly_idx[4:0]};
                addr_q_calc  = {bfly_idx[6:5], 1'b1, bfly_idx[4:0]};
                tw_addr_calc = {bfly_idx[4:0], 2'd0};
            end
            3'd6: begin
                addr_p_calc  = {bfly_idx[6], 1'b0, bfly_idx[5:0]};
                addr_q_calc  = {bfly_idx[6], 1'b1, bfly_idx[5:0]};
                tw_addr_calc = {bfly_idx[5:0], 1'd0};
            end
            3'd7: begin
                addr_p_calc  = {1'b0, bfly_idx[6:0]};
                addr_q_calc  = {1'b1, bfly_idx[6:0]};
                tw_addr_calc = bfly_idx[6:0];
            end
        endcase
    end

    // ======================================================================
    // Butterfly computation pipeline
    // ======================================================================

    // Latched values from registered RAM reads
    reg signed [15:0] a_re, a_im;
    reg signed [15:0] b_re, b_im;
    reg signed [15:0] tw_cos_r, tw_sin_r;
    reg [7:0] addr_p_r, addr_q_r;

    // Complex twiddle multiply: W * B
    // W = cos - j*sin, so W*B = (cos*Bre + sin*Bim) + j(cos*Bim - sin*Bre)
    wire signed [31:0] tw_x_re = tw_cos_r * b_re + tw_sin_r * b_im;
    wire signed [31:0] tw_x_im = tw_cos_r * b_im - tw_sin_r * b_re;

    // Scale twiddle product back from Q1.14 (arithmetic right shift by 14)
    wire signed [17:0] t_re = tw_x_re[31:14];
    wire signed [17:0] t_im = tw_x_im[31:14];

    // Butterfly results with 1/2 scaling per stage
    wire signed [17:0] a_re_ext = {{2{a_re[15]}}, a_re};
    wire signed [17:0] a_im_ext = {{2{a_im[15]}}, a_im};

    wire signed [17:0] sum_re = a_re_ext + t_re;
    wire signed [17:0] sum_im = a_im_ext + t_im;
    wire signed [17:0] dif_re = a_re_ext - t_re;
    wire signed [17:0] dif_im = a_im_ext - t_im;

    // Arithmetic right shift by 1, truncate to 16 bits
    wire [15:0] p_re_new = sum_re[16:1];
    wire [15:0] p_im_new = sum_im[16:1];
    wire [15:0] q_re_new = dif_re[16:1];
    wire [15:0] q_im_new = dif_im[16:1];

    // ======================================================================
    // Magnitude computation (from registered RAM reads during MAGNITUDE phase)
    // ======================================================================
    reg [7:0] mag_count;
    reg       mag_step;
    reg [7:0] mag_count_d;

    wire [15:0] abs_re = re_rdata_a[15] ? (~re_rdata_a + 16'd1) : re_rdata_a;
    wire [15:0] abs_im = im_rdata_a[15] ? (~im_rdata_a + 16'd1) : im_rdata_a;
    wire [15:0] mag_max = (abs_re > abs_im) ? abs_re : abs_im;
    wire [15:0] mag_min = (abs_re > abs_im) ? abs_im : abs_re;
    // Approximate magnitude: max + min/4 (within ~5% of true magnitude)
    wire [15:0] magnitude = mag_max + {2'b00, mag_min[15:2]};
    wire [15:0] scaled_mag = magnitude >> MAG_SHIFT;
    wire [8:0]  capped_mag = (scaled_mag > {7'd0, MAX_MAG}) ? MAX_MAG : scaled_mag[8:0];

    // ======================================================================
    // RAM port address/control mux (directly drives dual-port RAM signals)
    // ======================================================================
    always @(*) begin
        // Defaults: no writes, address 0
        re_addr_a  = 8'd0;  re_addr_b  = 8'd0;
        re_wdata_a = 16'd0; re_wdata_b = 16'd0;
        re_we_a    = 1'b0;  re_we_b    = 1'b0;
        im_addr_a  = 8'd0;  im_addr_b  = 8'd0;
        im_wdata_a = 16'd0; im_wdata_b = 16'd0;
        im_we_a    = 1'b0;  im_we_b    = 1'b0;
        tw_addr    = 7'd0;

        case (state)
            S_COLLECT: begin
                re_addr_a  = bit_reverse(sample_count);
                re_wdata_a = sample_in;
                re_we_a    = sample_valid;
                im_addr_a  = bit_reverse(sample_count);
                im_wdata_a = 16'd0;
                im_we_a    = sample_valid;
            end

            S_COMPUTE: begin
                tw_addr = tw_addr_calc;
                case (bfly_step)
                    2'd0: begin
                        // Read setup: present addresses for registered read
                        re_addr_a = addr_p_calc;
                        re_addr_b = addr_q_calc;
                        im_addr_a = addr_p_calc;
                        im_addr_b = addr_q_calc;
                    end
                    2'd1: begin
                        // Read data is now available in rdata registers
                        // (latching into a_re/b_re happens in state machine)
                    end
                    2'd2: begin
                        // Write butterfly results via both ports
                        re_addr_a  = addr_p_r;
                        re_addr_b  = addr_q_r;
                        re_wdata_a = p_re_new;
                        re_wdata_b = q_re_new;
                        re_we_a    = 1'b1;
                        re_we_b    = 1'b1;
                        im_addr_a  = addr_p_r;
                        im_addr_b  = addr_q_r;
                        im_wdata_a = p_im_new;
                        im_wdata_b = q_im_new;
                        im_we_a    = 1'b1;
                        im_we_b    = 1'b1;
                    end
                    default: ;
                endcase
            end

            S_MAGNITUDE: begin
                re_addr_a = mag_count;
                im_addr_a = mag_count;
            end

            default: ;
        endcase
    end

    // ======================================================================
    // Main state machine
    // ======================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state        <= S_COLLECT;
            sample_count <= 8'd0;
            bfly_stage   <= 3'd0;
            bfly_idx     <= 7'd0;
            bfly_step    <= 2'd0;
            mag_count    <= 8'd0;
            mag_step     <= 1'b0;
            mag_valid    <= 1'b0;
            mag_addr     <= 8'd0;
            mag_data     <= 9'd0;
        end else begin
            mag_valid <= 1'b0;  // Default: no output

            case (state)
                // ----------------------------------------------------------
                // COLLECT: Store 256 incoming samples at bit-reversed addresses
                // Writes are driven by the combinational mux above.
                // ----------------------------------------------------------
                S_COLLECT: begin
                    if (sample_valid) begin
                        if (sample_count == 8'd255) begin
                            sample_count <= 8'd0;
                            bfly_stage   <= 3'd0;
                            bfly_idx     <= 7'd0;
                            bfly_step    <= 2'd0;
                            state        <= S_COMPUTE;
                        end else begin
                            sample_count <= sample_count + 8'd1;
                        end
                    end
                end

                // ----------------------------------------------------------
                // COMPUTE: 8 stages x 128 butterflies x 3 cycles each
                // Step 0: present addresses (RAM reads on next posedge)
                // Step 1: latch registered read data + twiddle
                // Step 2: write butterfly results (via mux), advance
                // ----------------------------------------------------------
                S_COMPUTE: begin
                    case (bfly_step)
                        2'd0: begin
                            // Addresses driven by mux; latch for write-back
                            addr_p_r  <= addr_p_calc;
                            addr_q_r  <= addr_q_calc;
                            bfly_step <= 2'd1;
                        end
                        2'd1: begin
                            // Registered reads are now valid; latch into butterfly regs
                            a_re     <= $signed(re_rdata_a);
                            a_im     <= $signed(im_rdata_a);
                            b_re     <= $signed(re_rdata_b);
                            b_im     <= $signed(im_rdata_b);
                            tw_cos_r <= $signed(tw_rdata[31:16]);
                            tw_sin_r <= $signed(tw_rdata[15:0]);
                            bfly_step <= 2'd2;
                        end
                        2'd2: begin
                            // Writes driven by mux; advance to next butterfly
                            bfly_step <= 2'd0;
                            if (bfly_idx == 7'd127) begin
                                bfly_idx <= 7'd0;
                                if (bfly_stage == 3'd7) begin
                                    mag_count <= 8'd0;
                                    mag_step  <= 1'b0;
                                    state     <= S_MAGNITUDE;
                                end else begin
                                    bfly_stage <= bfly_stage + 3'd1;
                                end
                            end else begin
                                bfly_idx <= bfly_idx + 7'd1;
                            end
                        end
                        default: bfly_step <= 2'd0;
                    endcase
                end

                // ----------------------------------------------------------
                // MAGNITUDE: Compute |FFT[k]| for each bin, output to display
                // Step 0: present address (RAM read on next posedge)
                // Step 1: registered data valid → compute + output magnitude
                // ----------------------------------------------------------
                S_MAGNITUDE: begin
                    case (mag_step)
                        1'b0: begin
                            // Address driven by mux; save index for output
                            mag_count_d <= mag_count;
                            mag_step    <= 1'b1;
                        end
                        1'b1: begin
                            // Registered reads valid → compute magnitude combinationally
                            mag_addr  <= mag_count_d;
                            mag_data  <= capped_mag;
                            mag_valid <= 1'b1;
                            mag_step  <= 1'b0;
                            if (mag_count == 8'd255) begin
                                mag_count <= 8'd0;
                                state     <= S_COLLECT;
                            end else begin
                                mag_count <= mag_count + 8'd1;
                            end
                        end
                    endcase
                end

                default: state <= S_COLLECT;
            endcase
        end
    end

endmodule
